This is my first push in Git

This is my second change inthis file 

