This file will only showsup in new branch.
