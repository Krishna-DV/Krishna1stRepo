This is my first push in Git
